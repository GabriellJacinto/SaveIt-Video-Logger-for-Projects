*Library xor's finFET

*XOR V1
.subckt xor_1_fet a b xor vccbloco vssbloco vdd ground 
Mp1 vccbloco na nodo1 vdd                pmos_rvt w=27.0n l=20n nfin=1
Mp2 nodo1 b xor vdd                      pmos_rvt w=27.0n l=20n nfin=1
Mp3 vccbloco a nodo2 vdd                 pmos_rvt w=27.0n l=20n nfin=1
Mp4 nodo2 nb xor vdd                     pmos_rvt w=27.0n l=20n nfin=1
Mn1 xor nb nodo3 ground                  nmos_rvt w=27.0n l=20n nfin=1
Mn2 nodo3 na vssbloco ground             nmos_rvt w=27.0n l=20n nfin=1
Mn3 xor b nodo4 ground                   nmos_rvt w=27.0n l=20n nfin=1
Mn4 nodo4 a vssbloco ground              nmos_rvt w=27.0n l=20n nfin=1
Mpinv_a vccbloco a na vdd                pmos_rvt w=27.0n l=20n nfin=1
Mninv_a na a vssbloco ground             nmos_rvt w=27.0n l=20n nfin=1   
Mpinv_b vccbloco b nb vdd                pmos_rvt w=27.0n l=20n nfin=1
Mninv_b nb b vssbloco ground             nmos_rvt w=27.0n l=20n nfin=1
.ends xor_1_fet


*XOR V5
.subckt xor_5_fet a b xor vccbloco vssbloco vdd ground 
Mp1 a b xor vdd               				pmos_rvt w=27.0n l=20n nfin=1
Mp2 na nb xor vdd            				pmos_rvt w=27.0n l=20n nfin=1
Mn1 a nb xor ground           				nmos_rvt w=27.0n l=20n nfin=1
Mn2 na b xor ground          				nmos_rvt w=27.0n l=20n nfin=1
Mpinv_a vccbloco a na vdd          			pmos_rvt w=27.0n l=20n nfin=1
Mninv_a na a vssbloco ground    			nmos_rvt w=27.0n l=20n nfin=1  
Mpinv_b vccbloco b nb vdd          			pmos_rvt w=27.0n l=20n nfin=1
Mninv_b nb b vssbloco ground   				nmos_rvt w=27.0n l=20n nfin=1   
.ends xor_5_fet


*XOR V8
.subckt xor_8_fet a b xor vccbloco vssbloco vdd ground 
Mp1 vccbloco b nodo1 vdd            		pmos_rvt w=27.0n l=20n nfin=1
Mp2 a b xor vdd               				pmos_rvt w=27.0n l=20n nfin=1
Mp3 b a xor vdd               				pmos_rvt w=27.0n l=20n nfin=1
Mn1 nodo1 b vssbloco ground   				nmos_rvt w=27.0n l=20n nfin=1   
Mn2 a nodo1 xor ground   					nmos_rvt w=27.0n l=20n nfin=1   
Mn3 nodo1 a xor ground   					nmos_rvt w=27.0n l=20n nfin=1   
.ends xor_8_fet

*SOMADORES
.subckt cout_fet a cin h h_not cout vccbloco vssbloco vdd ground 
Mp1 cin h_not cout vdd            			pmos_rvt w=27.0n l=20n nfin=1
Mp2 a h cout vdd               				pmos_rvt w=27.0n l=20n nfin=1
Mn1 cin h cout ground   					nmos_rvt w=27.0n l=20n nfin=1  
Mn2 a h_not cout ground   					nmos_rvt w=27.0n l=20n nfin=1   
Mp3 vccbloco h h_not vdd            		pmos_rvt w=27.0n l=20n nfin=1
Mn3 h_not h vssbloco ground					nmos_rvt w=27.0n l=20n nfin=1   
.ends cout_fet


*-----------------------------------------------------------------------------
* Somador Mirror
*-----------------------------------------------------------------------------
.subckt mirror inCin inA inB Cout S vccbloco vssbloco vdd ground 

	Mp1 vccbloco inA a vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp2 a inB f vdd 							pmos_rvt w=27.0n l=20n nfin=1
	Mp3 vccbloco inA b vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp4 b inCin f vdd 							pmos_rvt w=27.0n l=20n nfin=1
	Mp5 vccbloco inB b vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp6 vccbloco inCin c vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp7 vccbloco inA c vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp8 vccbloco inB c vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp9 c f g vdd 								pmos_rvt w=27.0n l=20n nfin=1
	Mp10 vccbloco inA d vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp11 d inB e vdd 							pmos_rvt w=27.0n l=20n nfin=1
	Mp12 e inCin g vdd 							pmos_rvt w=27.0n l=20n nfin=1

	Mn1 f inB h ground 							nmos_rvt w=27.0n l=20n nfin=1 
	Mn2 h inA vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1 
	Mn3 i inA vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1 
	Mn4 f inCin i ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn5 i inB vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1
	Mn6 g f j ground 							nmos_rvt w=27.0n l=20n nfin=1
	Mn7 j inCin vssbloco ground 				nmos_rvt w=27.0n l=20n nfin=1
	Mn8 j inA vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1
	Mn9 j inB vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1
	Mn10 g inCin k ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn11 k inB l ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn12 l inA vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1

	*inversores
	Mp13 vccbloco g S vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mn13 S g vssbloco ground 					nmos_rvt w=27.0n l=20n nfin=1
	Mp14 vccbloco f Cout vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mn14 Cout f vssbloco ground 				nmos_rvt w=27.0n l=20n nfin=1

.ends

*-----------------------------------------------------------------------------
* Somador TGA
*-----------------------------------------------------------------------------
.subckt TGA inCin inA inB Cout S vccbloco vssbloco vdd ground 

	Mp1 vccbloco inB a vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp2 inA inB b vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp3 vccbloco inA c vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp4 c a b vdd 							pmos_rvt w=27.0n l=20n nfin=1
	Mp5 vccbloco inCin d vdd 				pmos_rvt w=27.0n l=20n nfin=1
	Mp6 inCin b S vdd 						pmos_rvt w=27.0n l=20n nfin=1
	Mp7 d e S vdd 							pmos_rvt w=27.0n l=20n nfin=1
	Mp8 vccbloco b e vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp9 inCin e Cout vdd 					pmos_rvt w=27.0n l=20n nfin=1
	Mp10 inA b Cout vdd 					pmos_rvt w=27.0n l=20n nfin=1

	Mn1 a inB vssbloco ground 				nmos_rvt w=27.0n l=20n nfin=1
	Mn2 inA a b ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn3 c inA vssbloco ground 				nmos_rvt w=27.0n l=20n nfin=1
	Mn4 c inB b ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn5 d inCin vssbloco ground 			nmos_rvt w=27.0n l=20n nfin=1
	Mn6 inCin e S ground 					nmos_rvt w=27.0n l=20n nfin=1
	Mn7 d b S ground 						nmos_rvt w=27.0n l=20n nfin=1
	Mn8 e b vssbloco ground 				nmos_rvt w=27.0n l=20n nfin=1
	Mn9 inCin b Cout ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn10 inA e Cout ground					nmos_rvt w=27.0n l=20n nfin=1
.ends

*----------------------------------------------
* Full adder TFA
*----------------------------------------------
.subckt TFA in_cin in_a in_b cout sum vccbloco vssbloco vdd ground 

	Mp1 vccbloco in_b p1_n1 vdd         	    pmos_rvt w=27.0n l=20n nfin=1
	Mp2 in_a in_b p3_p5 vdd        		        pmos_rvt w=27.0n l=20n nfin=1
	Mp3 in_b in_a p3_p5 vdd      	        	pmos_rvt w=27.0n l=20n nfin=1
	Mp4 in_cin p3_p5 sum vdd                	pmos_rvt w=27.0n l=20n nfin=1
	Mp5 p3_p5 in_cin sum vdd              		pmos_rvt w=27.0n l=20n nfin=1
	Mp6 vccbloco p3_p5 p6_n6 vdd                pmos_rvt w=27.0n l=20n nfin=1
	Mp7 in_cin p6_n6 cout vdd           	    pmos_rvt w=27.0n l=20n nfin=1
	Mp8 in_a p3_p5 cout vdd             	    pmos_rvt w=27.0n l=20n nfin=1

	Mn1 p1_n1 in_b vssbloco ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn2 in_a p1_n1 p3_p5 ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn3 p1_n1 in_a p3_p5 ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn4 in_cin p6_n6 sum ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn5 p6_n6 in_cin sum ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn6 p6_n6 p3_p5 vssbloco ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn7 in_cin p3_p5 cout ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn8 in_a p6_n6 cout ground					nmos_rvt w=27.0n l=20n nfin=1

.ends

*----------------------------------------------
* Full adder Hybrid
*----------------------------------------------
.subckt hybrid in_cin in_a in_b cout sum vccbloco vssbloco vdd ground 

	Mp1 in_a in_b p1_p2 vdd              	  	pmos_rvt w=27.0n l=20n nfin=1
	Mp2 p1_p2 in_a in_b vdd                		pmos_rvt w=27.0n l=20n nfin=1
	Mp3 vccbloco p1_p2 n1_p3 vdd                pmos_rvt w=27.0n l=20n nfin=1
	Mp4 vccbloco in_a p4_p5 vdd                	pmos_rvt w=27.0n l=20n nfin=1
	Mp5 p4_p5 in_b n1_p3 vdd                	pmos_rvt w=27.0n l=20n nfin=1
	Mp6 vccbloco in_cin p6_p7 vdd               pmos_rvt w=27.0n l=20n nfin=1
	Mp7 p6_p7 n1_p3 p7_n6 vdd             	    pmos_rvt w=27.0n l=20n nfin=1
	Mp8 vccbloco in_b p8_p9 vdd                 pmos_rvt w=27.0n l=20n nfin=1
	Mp9 p8_p9 in_a p7_n6 vdd                	pmos_rvt w=27.0n l=20n nfin=1
	Mp10 n10_n11 n1_p3 in_cin vdd               pmos_rvt w=27.0n l=20n nfin=1
	Mp11 n10_n11 in_cin n1_p3 vdd               pmos_rvt w=27.0n l=20n nfin=1
	
	Mn1 in_a in_b n1_p3 ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn2 n1_p3 in_a in_b ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn3 p1_p2 n1_p3 vssbloco ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn4 p1_p2 in_b n4_n5 ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn5 n4_n5 in_a vssbloco ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn6 p7_n6 p1_p2 n6_n7 ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn7 n6_n7 in_cin vssbloco ground			nmos_rvt w=27.0n l=20n nfin=1
	Mn8 p7_n6 in_a n8_n9 ground					nmos_rvt w=27.0n l=20n nfin=1
	Mn9 n8_n9 in_b vssbloco ground				nmos_rvt w=27.0n l=20n nfin=1
	Mn10 in_cin p1_p2 n10_n11 ground			nmos_rvt w=27.0n l=20n nfin=1
	Mn11 p1_p2 in_cin n10_n11 ground			nmos_rvt w=27.0n l=20n nfin=1

	*inversores
	Mp12 vccbloco n10_n11 sum vdd 				pmos_rvt w=27.0n l=20n nfin=1
	Mn12 sum n10_n11 vssbloco ground 			nmos_rvt w=27.0n l=20n nfin=1
	Mp13 vccbloco p7_n6 cout vdd 				pmos_rvt w=27.0n l=20n nfin=1
	Mn13 cout p7_n6 vssbloco ground 			nmos_rvt w=27.0n l=20n nfin=1
	
.ends

*Fim do Arquivo SPICE
*.end
