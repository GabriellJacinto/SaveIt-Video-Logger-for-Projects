*FA_VxVx.cir

*Modelo do transistor
***** PARAMETROS
		.include "7nm_FF.pm"
		.include LIBRARY_FinFET_traditional.cir
        .param supply = 0.35V
        .param ground_valor = 0
        .temp 0 25 50 75 100 125 
******
.global vdd gnd ground wfn wfp
******************************************************************
		.include fontes_SOMA.cir
		.include ondas_SOMA.cir
		.include inversores_in_out_SOMA.cir
		
*****INSTANCIA��O DO SUBCKT(SOMADORES)
		X1 cin1 a1 b1 cout sum vccbloco vssbloco vdd ground mirror          
******
*****TIPO DE SIMULA��O
		.tran 1p 144n 
******	
		.include atrasos_SOMA.cir
		.include energia_SOMA.cir
		.include potencia_SOMA.cir
******************************************************************

*Fim do Arquivo SPICE
.end


